module i2s #(
    parameter SYS_CLK     = 50_000_000,  // ϵͳ�ο�ʱ��
    parameter SAMPLE_RATE = 48_000,      // I2S������
    parameter DEPTH       = 16           // ����λ������
)(
    input                    clk_50m,     // ����ο�ʱ��
    input                    rst_n,       // �͵�ƽ��λ
    input                    ADC_DAT,     // ������ƵADC��������
    output                   BCLK,        // ���i2s��Ƶʱ��
    output                   ADC_LRC,     // ���ADC���������ź�
    output                   DAC_LRC,     // ���DAC���������ź�
    output [31:0]            o_rx_data    // ����ADC���ݣ�����32λ�ӿڲ��䣩
);

    // BLCK����ź�
    wire p_bclk;
    wire n_bclk;

    // i2sʱ������ģ�飨��������WM8731Ϊ�ӻ�
    timing_gen #(
        .SYS_CLK             (SYS_CLK)     ,
        .SAMPLE_RATE         (SAMPLE_RATE) ,
        .DEPTH               (DEPTH)
    ) u_timing_gen (
        .clk_50m             (clk_50m)     ,
        .rst_n               (rst_n)       ,
        .BCLK                (BCLK)        ,
        .ADC_LRC             (ADC_LRC)     ,
        .DAC_LRC             (DAC_LRC)     ,
        .p_bclk              (p_bclk)      ,
        .n_bclk              (n_bclk)
    );

    // ��Ƶ���մ�ת��
    rx #(
        .DEPTH (DEPTH)
    ) u_rx (
        .clk_50m             (clk_50m)     ,
        .rst_n               (rst_n)       ,
        .ADC_LRC             (ADC_LRC)     ,
        .ADC_DAT             (ADC_DAT)     ,
        .i_p_bclk            (p_bclk)      ,
        .i_n_bclk            (n_bclk)      ,
        .o_rx_data           (o_rx_data)
    );

endmodule
