module top_codec( 
    input  clk_50m                      ,    // ����ο�ʱ��   
    input  rst_n                        ,    // �͵�ƽ��λ     
    input  ADC_DAT                      ,    // ������ƵADC��������   
    output BCLK                         ,    // ���i2s��Ƶʱ��       
    output ADC_LRC                      ,    // ���ADC���������ź�       
    output DAC_LRC                      ,    // ���DAC���������ź�       
    output DAC_DAT                      ,    // �����ƵDAC�������ݣ�����ԭ�˿ڣ�δ������
    output I2C_SCLK                     ,    // i2c���� SCL
    inout  I2C_SDAT                          // i2c���� SDA
);

    // ���н�������
    wire [31:0] o_rx_data;

    i2s #(
        .SYS_CLK      (50_000_000)      ,
        .SAMPLE_RATE  (48_000)          ,
        .DEPTH        (16)
    ) u_i2s (
        .clk_50m      (clk_50m)         ,
        .rst_n        (rst_n)           ,
        .ADC_DAT      (ADC_DAT)         ,
        .BCLK         (BCLK)            ,
        .ADC_LRC      (ADC_LRC)         ,
        .DAC_LRC      (DAC_LRC)         ,
        .o_rx_data    (o_rx_data)
    );


    i2c u_i2c(
        .clk_50m      (clk_50m)         ,
        .rst_n        (rst_n)           ,
        .I2C_SCLK     (I2C_SCLK)        ,
        .I2C_SDAT     (I2C_SDAT)
    );


endmodule
