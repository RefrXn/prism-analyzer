module i2c(
    input        clk_50m                ,    // ʱ���ź�
    input        rst_n                  ,    // ��λ�ź�
    
	output       i2c_ack                ,    // I2CӦ���־ 0:Ӧ�� 1:δӦ��
    output       I2C_SCLK               ,    // wm8731��SCLʱ��
    inout        I2C_SDAT                    // wm8731��SDA�ź�
);

    //parameter define
    parameter   SLAVE_ADDR = 7'h1a         ;    // ������ַ
    parameter   WL         = 6'd32         ;    // word length��Ƶ�ֳ���������
    parameter   BIT_CTRL   = 1'b0          ;    // �ֵ�ַλ���Ʋ���(16b/8b)
    parameter   CLK_FREQ   = 30'd50_000_000;    // i2c_driģ�������ʱ��Ƶ��(CLK_FREQ)
    parameter   I2C_FREQ   = 18'd250_000   ;    // I2C��SCLʱ��Ƶ��
    
    //wire define
    wire        clk_i2c   ;                     // i2c�Ĳ���ʱ��
    wire        i2c_exec  ;                     // i2c��������
    wire        i2c_done  ;                     // i2c����������־
    wire        cfg_done  ;                     // wm8731������ɱ�־
    wire [15:0] reg_data  ;                     // wm8731��Ҫ���õļĴ�������ַ�����ݣ�
    
    
    
    //����wm8731�ļĴ���
    i2c_reg_cfg u_i2c_reg_cfg(  
        .clk_i2c        (clk_i2c        ),       // i2c_reg_cfg����ʱ��
        .rst_n          (rst_n          ),       // ��λ�ź�
      
        .i2c_exec       (i2c_exec       ),       // I2C����ִ���ź�
        .i2c_data       (reg_data       ),       // �Ĵ������ݣ�7λ��ַ+9λ���ݣ�
        
        .i2c_done       (i2c_done       ),       // I2Cһ�β�����ɵı�־�ź�            
        .cfg_done       (cfg_done       )        // wm8731�������
    );
    
    //����IICЭ��
    i2c_dri #(
        .SLAVE_ADDR     (SLAVE_ADDR),            // slave address�ӻ���ַ���Ŵ˴������������
        .CLK_FREQ       (CLK_FREQ       ),       // i2c_driģ�������ʱ��Ƶ��(CLK_FREQ)
        .I2C_FREQ       (I2C_FREQ       )        // I2C��SCLʱ��Ƶ��
    ) u_i2c_dri(  
        .clk_50m        (clk_50m        ),       // i2c_driģ�������ʱ��(CLK_FREQ)
        .rst_n          (rst_n          ),       // ��λ�ź�
      
        .i2c_exec       (i2c_exec       ),       // I2C����ִ���ź�
        .bit_ctrl       (BIT_CTRL       ),       // ������ַλ����(16b/8b)
        .i2c_rh_wl      (1'b0           ),       // I2C��д�����ź�
        .i2c_addr       (reg_data[15:8] ),       // I2C�����ֵ�ַ
        .i2c_data_w     (reg_data[ 7:0] ),       // I2CҪд������
          
        .i2c_done       (i2c_done       ),       // I 2Cһ�β������
        .i2c_ack        (i2c_ack        ),       // I2CӦ���־ 0:Ӧ�� 1:δӦ��
          
        .scl            (I2C_SCLK       ),       // I2C��SCLʱ���ź�
        .sda            (I2C_SDAT       ),       // I2C��SDA�ź�
        .dri_clk        (clk_i2c        )        // I2C����ʱ��
    );
    
endmodule 