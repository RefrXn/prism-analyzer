module band_accum #(
    parameter integer FFT_LEN   = 1024,  // FFT ������������ 2 ���ݣ�
    parameter integer BANDS     = 32,    // ���Ƶ����
    parameter integer IN_WIDTH  = 24,    // �������λ��
    parameter integer OUT_WIDTH = 16     // �������λ��
) (
    input  wire                     clk_50m,
    input  wire                     rst_n,

    // ���룺ÿ֡ N ��ķ��ȣ��� FFT ������룩��ֻͳ�� [0 .. N/2-1] �� N/2 ��
    // NOTE: FFT ����� DC ������ tdata[0] ��������
    input  wire                     s_axis_tvalid,
    output wire                     s_axis_tready,
    input  wire [IN_WIDTH-1:0]      s_axis_tdata,
    input  wire                     s_axis_tlast,

    // �����ÿ֡���� BANDS ��ֵ��������ͺ��λ�������һ���� tlast
    output reg                      m_axis_tvalid,
    input  wire                     m_axis_tready,
    output      [OUT_WIDTH-1:0]     m_axis_tdata,
    output reg                      m_axis_tlast
);

    // ===============================================================
    // 1) ������ֲ�����
    // ===============================================================
    localparam integer HALF_N       = FFT_LEN / 2;
    localparam integer BAND_SAMPLES = HALF_N / BANDS;

    // ===============================================================
    // 2) �Ĵ�������
    // ===============================================================
    reg [$clog2(BAND_SAMPLES):0]            band_sample_idx;  // ��ǰ band �ڲ���������
    reg [$clog2(BANDS):0]                   band_idx;         // ��ǰ�ۼӵ��ڼ��� band
    reg [IN_WIDTH+$clog2(BAND_SAMPLES)-1:0] acc, acc_r;       // �ۼ���
    reg                                     frame_done;

    // �����λӳ��
    assign m_axis_tdata = acc_r[IN_WIDTH+$clog2(BAND_SAMPLES)-1-:OUT_WIDTH];

    // ���� ready ����
    assign s_axis_tready = (!m_axis_tvalid) || m_axis_tready;

    // ===============================================================
    // 3) ��ʱ���߼�
    // ===============================================================
    always @(posedge clk_50m) begin
        if (!rst_n) begin
            band_sample_idx <= 0;
            band_idx        <= 0;
            acc             <= 0;
            acc_r           <= 0;
            m_axis_tvalid   <= 0;
            m_axis_tlast    <= 0;
            frame_done      <= 0;
        end
        else begin
            // -------------------------------------------------------
            // �������ֺ��� valid
            // -------------------------------------------------------
            if (m_axis_tvalid && m_axis_tready) begin
                m_axis_tvalid <= 1'b0;
                m_axis_tlast  <= 1'b0;
            end

            // -------------------------------------------------------
            // ���봦��
            // -------------------------------------------------------
            if (s_axis_tvalid && s_axis_tready) begin
                if (!frame_done) begin
                    // =======================
                    // ��ǰ band �����ۼ�
                    // =======================
                    if (band_sample_idx == BAND_SAMPLES - 1) begin
                        // ��ǰ band �ۼ���ɣ�������
                        acc             <= 'b0;
                        acc_r           <= acc + s_axis_tdata;
                        m_axis_tvalid   <= 1'b1;
                        m_axis_tlast    <= (band_idx == BANDS - 1) ? 1'b1 : 1'b0;
                        band_sample_idx <= 0;
                        band_idx        <= band_idx + 1;
                        frame_done      <= (band_idx == BANDS - 1) ? 1'b1 : 1'b0;
                    end
                    else begin
                        // �����ۼӵ�ǰ band
                        acc             <= (band_sample_idx == 0 && band_idx == 0) ?
                                            s_axis_tdata : acc + s_axis_tdata;
                        band_sample_idx <= band_sample_idx + 1;
                    end
                end
                else begin
                    // =======================
                    // ֡������λ״̬
                    // =======================
                    if (s_axis_tlast) begin
                        band_sample_idx <= 'b0;
                        band_idx        <= 'b0;
                        acc             <= 'b0;
                        frame_done      <= 1'b0;
                    end
                end
            end
        end
    end

endmodule
