`timescale 1ns / 1ps
module ws2812_dri (
    input              clk_50m      ,     // 50MHz ʱ������
    input              rst_n        ,     // ��λ�źţ�����Ч��
    input  wire        start        ,     // ֡��ʼ����һ�ģ�
    input  wire        valid        ,     // ������Ч�����������ڼ�ÿ�����ش�һ�� done_bit��
    input  wire [23:0] din          ,     // GRB ��������
    output reg         dout         ,     // WS2812 ������
    output reg         done_bit     ,     // �������ش�����ɣ���һ�ģ�
    output reg         done_dz            // ȫ��������ɣ���λʱ�������һ�ģ�
);

    // WS2812B ʱ����� (50MHz������20ns)
    parameter T0H = 17              ;     // 0 �ߵ�ƽ ~340ns
    parameter T1H = 45              ;     // 1 �ߵ�ƽ ~900ns
    parameter T0L = 35              ;     // 0 �͵�ƽ ~700ns
    parameter T1L = 27              ;     // 1 �͵�ƽ ~540ns
    parameter RESET_CYCLES = 14000  ;     // >280us ��λ

    reg [13:0] cnt                   ;     // ���ڼ���
    reg [ 4:0] cnt_bit               ;     // 24bit����
    reg [ 8:0] cnt_bety              ;     // 256�ŵƼ���
    reg [23:0] data_reg              ;     // ��ǰ�������ݼĴ�
    reg [ 6:0] cur_state, next_state ;

    // FSM ״̬����
    localparam  IDLE = 7'b0000001    , 
                START = 7'b0000010   , 
                DATA0 = 7'b0000100   , 
                DATA1 = 7'b0001000   , 
                ACK = 7'b0010000     , 
                STOP = 7'b0100000    , 
                RES = 7'b1000000     ;

    // ״̬��ʱ��
    always @(posedge clk_50m or negedge rst_n) begin
        if (!rst_n) cur_state <= IDLE;
        else cur_state <= next_state;
    end

    // ״̬�����
    always @(*) begin
        if (!rst_n) next_state = IDLE;
        else begin
            case (cur_state)
                IDLE  : next_state = (start || valid) ? START : IDLE;
                START : next_state = (data_reg[23-cnt_bit]==1'b0) ? DATA0 : DATA1;
                DATA0 : next_state = (cnt==T0H+T0L-1) ? ACK : DATA0;
                DATA1 : next_state = (cnt==T1H+T1L-1) ? ACK : DATA1;
                ACK   : next_state = (cnt_bit==5'd23) ? STOP : START;
                STOP  : next_state = (cnt_bety==9'd255) ? RES : IDLE;
                RES   : next_state = (cnt==RESET_CYCLES-1) ? IDLE : RES;
                default: next_state = IDLE;
            endcase
        end
    end

    // ��������
    always @(posedge clk_50m or negedge rst_n) begin
        if (!rst_n) begin
            data_reg <= 24'd0;
            cnt      <= 14'd0;
            cnt_bit  <= 5'd0;
            cnt_bety <= 9'd0;
            dout     <= 1'b0;
            done_bit <= 1'b0;
            done_dz  <= 1'b0;
        end else begin
            case (cur_state)
                IDLE: begin
                    data_reg <= din;  // �ڽ��� START ǰץȡ������
                    cnt_bety <= start ? 'b0 : cnt_bety;
                    cnt      <= 14'd0;
                    cnt_bit  <= 5'd0;
                    dout     <= 1'b0;
                    done_bit <= 1'b0;
                    done_dz  <= 1'b0;
                end

                START: begin
                    cnt      <= 14'd0;
                    dout     <= 1'b0;
                    done_bit <= 1'b0;
                    done_dz  <= 1'b0;
                end

                DATA0: begin
                    cnt      <= (cnt == T0H + T0L - 1) ? 14'd0 : cnt + 14'd1;
                    dout     <= (cnt < T0H);
                    done_bit <= 1'b0;
                    done_dz  <= 1'b0;
                end

                DATA1: begin
                    cnt      <= (cnt == T1H + T1L - 1) ? 14'd0 : cnt + 14'd1;
                    dout     <= (cnt < T1H);
                    done_bit <= 1'b0;
                    done_dz  <= 1'b0;
                end

                ACK: begin
                    cnt      <= 14'd0;
                    dout     <= 1'b0;
                    cnt_bit  <= (cnt_bit == 5'd23) ? 5'd0 : (cnt_bit + 5'd1);
                    done_dz  <= 1'b0;
                    done_bit <= 1'b0;
                end

                STOP: begin
                    cnt      <= 14'd0;
                    cnt_bety <= (cnt_bety == 9'd255) ? 9'd0 : (cnt_bety + 9'd1);
                    cnt_bit  <= 5'd0;
                    dout     <= 1'b0;
                    done_bit <= 1'b1;  // ��֪����"��ǰ���ط������"
                    done_dz  <= 1'b0;
                end

                RES: begin
                    if (cnt == RESET_CYCLES - 1) begin
                        cnt     <= 14'd0;
                        done_dz <= 1'b1;  // ȫ֡��λ���
                    end else begin
                        cnt     <= cnt + 14'd1;
                        done_dz <= 1'b0;
                    end
                    cnt_bety <= 9'd0;
                    cnt_bit  <= 5'd0;
                    dout     <= 1'b0;
                    done_bit <= 1'b0;
                end

                default: begin
                    data_reg <= 24'd0;
                    cnt      <= 14'd0;
                    cnt_bety <= 9'd0;
                    cnt_bit  <= 5'd0;
                    dout     <= 1'b0;
                    done_bit <= 1'b0;
                    done_dz  <= 1'b0;
                end
            endcase
        end
    end

endmodule
