// ===============================================================
// - ����: 16-bit PCM ���� (pcm_in_valid, pcm_in_sample)
// - ���: 32 ·Ƶ��ֵ (ͨ�� spectrum_out_ram ���ڵ���)
// ===============================================================
module top_fft #(
    parameter                             PCM_WIDTH           = 16       ,
    parameter                             FFT_LEN             = 1024     ,      
    parameter                             FFT_RE_IM_WIDTH     = 16       ,      // FFT IP ��ʵ��λ��(ÿ·)
    parameter                             MAG_WIDTH           = 16       ,      // ����λ���ڲ���
    parameter                             BANDS               = 32       ,      // Ŀ��Ƶ����
    parameter                             PEAK_HOLD_FRAMES    = 3                         // ��ֵ����֡��
)(
    input  wire                            clk_50m            ,
    input  wire                            rst_n              ,
        
    // PCM ���루����ʱ��48kHz����Чʱ����1�ļ��ɣ�
    input  wire                            pcm_in_valid       ,
    input  wire signed [PCM_WIDTH-1:0]     pcm_in_sample      ,

    // Ƶ�׶��ڣ������� WS2812 ģ�����ԣ�
    input  wire [clog2_fn(BANDS)-1:0]      spec_rd_addr       ,
    input  wire                            spec_rd_en         ,
    output wire [15:0]                     spec_rd_data       ,      // ѹ������� 16bit
    output wire                            spec_frame_stb     ,      // ÿ֡�������� 32 band����һ��
    output wire                            spec_rd_data_valid
);

    // 1) PCM -> AXIS (complex), ֡���
    wire                                   s_axis_tvalid      ;
    wire                                   s_axis_tready      ;
    wire [2*FFT_RE_IM_WIDTH-1:0]           s_axis_tdata       ;      // {Re, Im}
    wire                                   s_axis_tlast       ;

    frame_packer #(
        .PCM_WIDTH                         (PCM_WIDTH       )  ,
        .FFT_LEN                           (FFT_LEN         )  ,
        .FFT_RE_IM_WIDTH                   (FFT_RE_IM_WIDTH )
    ) u_frame_packer (
        .clk_50m                           (clk_50m         )  ,
        .rst_n                             (rst_n           )  ,
        .pcm_in_valid                      (pcm_in_valid    )  ,
        .pcm_in_sample                     (pcm_in_sample   )  ,
        .s_axis_tvalid                     (s_axis_tvalid   )  ,
        .s_axis_tready                     (s_axis_tready   )  ,
        .s_axis_tdata                      (s_axis_tdata    )  ,
        .s_axis_tlast                      (s_axis_tlast    )
    );


    // 2) FFT IP ��װ (AXIS in/out)
    wire                                   m_axis_tvalid       ;
    wire                                   m_axis_tready       ;
    wire [2*FFT_RE_IM_WIDTH-1:0]           m_axis_tdata        ;      // {Re, Im}
    wire                                   m_axis_tlast        ;

    fft_wrapper #(
        .FFT_LEN                           (FFT_LEN         )  ,
        .FFT_RE_IM_WIDTH                   (FFT_RE_IM_WIDTH )
    ) u_fft_wrapper (
        // Clock & Reset
        .clk_50m                           (clk_50m         )  ,
        .rst_n                             (rst_n           )  ,
        // S_AXIS (input)
        .s_axis_tvalid                     (s_axis_tvalid   )  ,
        .s_axis_tready                     (s_axis_tready   )  ,
        .s_axis_tdata                      (s_axis_tdata    )  ,
        .s_axis_tlast                      (s_axis_tlast    )  ,
        // M_AXIS (output)
        .m_axis_tvalid                     (m_axis_tvalid   )  ,
        .m_axis_tready                     (m_axis_tready   )  ,
        .m_axis_tdata                      (m_axis_tdata    )  ,
        .m_axis_tlast                      (m_axis_tlast    )
    );


    // 3) ���� -> ���ȣ����ƣ�
    wire                                   mag_tvalid          ;
    wire                                   mag_tready          ;
    wire [MAG_WIDTH-1:0]                   mag_tdata           ;
    wire                                   mag_tlast           ;
    
    assign spec_frame_stb = mag_tlast; // ������һ������ʱupdate

    complex_to_mag #(
        .RE_IM_WIDTH                       (FFT_RE_IM_WIDTH )  ,
        .MAG_WIDTH                         (MAG_WIDTH       )
    ) u_complex_to_mag (
        // Clock & Reset
        .clk_50m                           (clk_50m         )  ,
        .rst_n                             (rst_n           )  ,
        // S_AXIS (input)
        .s_axis_tvalid                     (m_axis_tvalid   )  ,
        .s_axis_tready                     (m_axis_tready   )  ,
        .s_axis_tdata                      (m_axis_tdata    )  ,  // {Re, Im}
        .s_axis_tlast                      (m_axis_tlast    )  ,
        // M_AXIS (output)
        .m_axis_tvalid                     (mag_tvalid      )  ,
        .m_axis_tready                     (mag_tready      )  ,
        .m_axis_tdata                      (mag_tdata       )  ,
        .m_axis_tlast                      (mag_tlast       )
    );
    
    
    // 4) Ƶ����� (N/2 -> 32 bands), ����ƽ��
    //    �˴����� DC(0) �� Nyquist(N/2)
    wire                                   band_tvalid         ;
    wire                                   band_tready         ;
    wire [15:0]                            band_tdata          ;   // �Ƚس�16λ����������ѹ��/��ֵ����
    wire                                   band_tlast          ;   // ÿ���һ�� band����һ�� valid�����һ�� band �� tlast������һ��band��һ��

    band_accum #(
        .FFT_LEN                           (FFT_LEN         )  ,
        .BANDS                             (BANDS           )  ,
        .IN_WIDTH                          (MAG_WIDTH       )  ,
        .OUT_WIDTH                         (16              )
    ) u_band_accum (
        // Clock & Reset
        .clk_50m                           (clk_50m         )  ,
        .rst_n                             (rst_n           )  ,
        // S_AXIS (input)
        .s_axis_tvalid                     (mag_tvalid      )  ,
        .s_axis_tready                     (mag_tready      )  ,
        .s_axis_tdata                      (mag_tdata       )  ,
        .s_axis_tlast                      (mag_tlast       )  ,
        // M_AXIS (output)
        .m_axis_tvalid                     (band_tvalid     )  ,
        .m_axis_tready                     (band_tready     )  ,
        .m_axis_tdata                      (band_tdata      )  ,
        .m_axis_tlast                      (band_tlast      )
    );


    // 5) ��ֵ���� + ����ѹ����log2���ƣ�
    wire                                   comp_tready                   ;
    wire                                   comp_tvalid = band_tvalid     ;
    wire [15:0]                            comp_tdata = band_tdata       ;
    wire                                   comp_tlast = band_tlast       ;
    
    assign                                 band_tready = comp_tready     ;


    // 6) д�� 32��16 RAM�����ⲿ��
    band_buffer #(
        .BANDS                             (BANDS           )  ,
        .DATA_WIDTH                        (16              )
    ) u_band_buffer (
        // Clock & Reset
        .clk_50m                           (clk_50m         )  ,
        .rst_n                             (rst_n           )  ,
    
        // д������ comp ����ÿ֡����д 0..BANDS-1
        .s_axis_tvalid                     (comp_tvalid     )  ,
        .s_axis_tready                     (comp_tready     )  ,
        .s_axis_tdata                      (comp_tdata      )  ,
        .s_axis_tlast                      (comp_tlast      )  ,
    
        // �����첽һ�ķ���
        .rd_addr                           (spec_rd_addr    )  ,
        .rd_en                             (spec_rd_en      )  ,
        .rd_data                           (spec_rd_data    )  ,
        .frame_stb                         (                )  ,  // ���ź��� FFT ��֡ʱ����������ã�Ӧ���� mag_tlast, ֮ǰ�ȹ���
        .rd_data_valid                     (spec_rd_data_valid)
    );

    
    // 7�����ƺ�����Ҳ������CORDIC���������ӳ�
    function   integer clog2_fn ;
        input  integer v        ;
               integer i        ;
        begin
            v = v - 1            ;
            for (i = 0; v > 0; i = i + 1)
                v = v >> 1       ;
            clog2_fn = i         ;
        end
    endfunction


endmodule
