module rx #(
    parameter DEPTH = 16                        // ÿ��������λ��
)(
    input  wire             clk_50m    ,        // ϵͳʱ�ӣ��� BCLK ͬ����
    input  wire             rst_n      ,        // �첽��λ���͵�ƽ��Ч
    input  wire             ADC_LRC    ,        // LRCLK����������ѡ���ź�
    input  wire             ADC_DAT    ,        // ���� ADC ��Ƶ����
    input  wire             i_p_bclk   ,        // BCLK ���ر�־
    input  wire             i_n_bclk   ,        // BCLK ���ر�־

    output reg  [DEPTH-1:0] o_rx_data  ,        // ��������յĲ�����Ƶ����
    output reg              o_rx_done           // �����һ֡������ɱ�־��1clk ��Ч��
);

    //============================================================
    // �ڲ��źŶ���
    //============================================================
    reg [7:0] rx_cnt;                           // bit λ������
    reg [DEPTH-1:0] r_rx_data;                  // ������λ�Ĵ���
    reg r_adc_rlc;                              // LRCLK �ӳټĴ���
    wire adc_rlc_edge;                          // LRCLK ��ת����ź�

    assign adc_rlc_edge = ADC_LRC ^ r_adc_rlc;  // ����ⷭת��

    //============================================================
    // LRCLK ���ؼ��
    //============================================================
    // ���� i_adc_rlc ��ǰһ�ģ����ڼ�����������л�ʱ��
    always @(posedge clk_50m) begin
        if (!rst_n)
            r_adc_rlc <= 1'b0;
        else if (i_n_bclk)
            r_adc_rlc <= ADC_LRC;
    end

    //============================================================
    // bit �����߼�
    //============================================================
    // ÿ֡����λ�� = SAMPLE_DEEP
    // LRCLK ��ת�����¼���
    always @(posedge clk_50m) begin
        if (!rst_n)
            rx_cnt <= 8'd0;
        else if (adc_rlc_edge)
            rx_cnt <= 8'd0;
        else if (rx_cnt < DEPTH + 8'd3 && i_p_bclk)
            rx_cnt <= rx_cnt + 8'd1;
    end

    //============================================================
    // ����������λ�Ĵ���
    //============================================================
    // �� BCLK ���ز�������Ĵ�������
    always @(posedge clk_50m) begin
        if (!rst_n)
            r_rx_data <= {DEPTH{1'b0}};
        else if (rx_cnt < DEPTH && i_p_bclk)
            r_rx_data <= {r_rx_data[DEPTH-2:0], ADC_DAT};
    end

    //============================================================
    // ��������Ĵ���
    //============================================================
    // ���������� SAMPLE_DEEP ʱ��������
    always @(posedge clk_50m) begin
        if (!rst_n)
            o_rx_data <= {DEPTH{1'b0}};
        else if (rx_cnt == DEPTH && i_p_bclk)
            o_rx_data <= r_rx_data;
    end

    //============================================================
    // ��������ź�
    //============================================================
    // o_rx_done ��ÿ֡���ս���ʱ����һ��ʱ������
    always @(posedge clk_50m) begin
        if (!rst_n)
            o_rx_done <= 1'b0;
        else if (rx_cnt == DEPTH && i_p_bclk)
            o_rx_done <= 1'b1;
        else
            o_rx_done <= 1'b0;
    end

endmodule
