module i2c_reg_cfg (
    input                clk_i2c  ,     // i2c_reg_cfg����ʱ��
    input                rst_n    ,     // ��λ�ź�
    input                i2c_done ,     // I2Cһ�β�����ɷ����ź�
    output  reg          i2c_exec ,     // I2C����ִ���ź�
    output  reg          cfg_done ,     // WM8978�������
    output  reg  [15:0]  i2c_data       // �Ĵ������ݣ�7λ��ַ+9λ���ݣ�
);

    localparam REG_NUM      = 5'd11;        // �ܹ���Ҫ���õļĴ�������
    localparam PHONE_LVOLUME = 7'd0;        // �������������������С������0~127��
    localparam PHONE_RVOLUME = 7'd120;        // �������������������С������0~127��
    
    
    
    //reg define
    reg    [7:0]  start_init_cnt;           // ��ʼ����ʱ������
    reg    [4:0]  init_reg_cnt  ;           // �Ĵ������ø���������
    
    //*****************************************************
    //**                    main code
    //*****************************************************
    
    //�ϵ��λ����ʱһ��ʱ��
    always @(posedge clk_i2c or negedge rst_n) begin
        if(!rst_n)
            start_init_cnt <= 8'd0;
        else if(start_init_cnt < 8'hff)
            start_init_cnt <= start_init_cnt + 1'b1;
    end
    
    //����I2C����
    always @(posedge clk_i2c or negedge rst_n) begin
        if(!rst_n)
            i2c_exec <= 1'b0;
        else if(init_reg_cnt == 5'd0 & start_init_cnt == 8'hfe)
            i2c_exec <= 1'b1;
        else if(i2c_done && init_reg_cnt < REG_NUM)
            i2c_exec <= 1'b1;
        else
            i2c_exec <= 1'b0;
    end
    
    //���üĴ�������
    always @(posedge clk_i2c or negedge rst_n) begin
        if(!rst_n)
            init_reg_cnt <= 5'd0;
        else if(i2c_exec)
            init_reg_cnt <= init_reg_cnt + 1'b1;
    end
    
    //�Ĵ�����������ź�
    always @(posedge clk_i2c or negedge rst_n) begin
        if(!rst_n)
            cfg_done <= 1'b0;
        else if(i2c_done & (init_reg_cnt == REG_NUM) )
            cfg_done <= 1'b1;
    end
    
    //����I2C�����ڼĴ�����ַ��������
    always @(posedge clk_i2c or negedge rst_n) begin
        if(!rst_n)
            i2c_data <= 16'b0;
        else begin
            case(init_reg_cnt)                    
                5'd0 : i2c_data <= {7'h0f ,9'b0};					// R15,��λ                    
                5'd1 : i2c_data <= {7'h00 ,9'b0_0001_0111};			// R0,δ�õ�                   
                5'd2 : i2c_data <= {7'h01 ,9'b0_0001_0111};			// R1,δ�õ�                 
                5'd3:  i2c_data <= {7'h02 ,{2'b01,PHONE_LVOLUME}};	// R2,��������������                   
                5'd4 : i2c_data <= {7'h03 ,{2'b01,PHONE_RVOLUME}};	// R3,��������������     
                5'd5 : i2c_data <= {7'h04 ,9'b0_0001_0100};         // R4,ʹ����˷磬�ر�mic����(������bypass),ȡ��mic���������
                5'd6 : i2c_data <= {7'h05 ,9'b0000_00110};			// R5,������Ƶ�������,�ر�adc����
                5'd7 : i2c_data <= {7'h06 ,9'b0_0000_0000};			// R6,power down
                5'd8 : i2c_data <= {7'h07 ,9'b0_0001_0010};			// R7,I2S,16bit,LRC(H)-->right ch,slave
                5'd9 : i2c_data <= {7'h08 ,9'b0_0000_0000};			// R8,ADC-->48K  DAC-->48K
                5'd10: i2c_data <= {7'h09 ,9'b0_0000_0001};			//ACTIVE
                default : ;
            endcase
        end
    end

endmodule 